`ifndef _incname_vh_
`define _incname_vh_


`endif //_incname_vh_
