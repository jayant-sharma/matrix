`define WIDTH 	16
`define MAT_SZ 	3
`define N	MAT_SZ

